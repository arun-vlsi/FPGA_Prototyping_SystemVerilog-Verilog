`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 16.10.2025 11:03:12
// Design Name: 
// Module Name: font_test_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module font_test_top
(
input wire clk, reset,
output wire hsync, vsync,
output wire [2:0] rgb
);

// signal declaration 
wire [9:0] pixel_x, pixel_y;
wire video_on, pixel_tick; 
reg [2:0] rgb_reg;
wire [2:0] rgb_next;

// body 
// instantiate vga sync circuit 
vga_sync vsync_unit(.clk(clk), .reset(reset), .hsync(hsync), .vsync(vsync),
                     .video_on(video_on), .p_tick(picel_tick),
                     .pixel_x(pixel_), .pixel_y(pixel_y));
 // font generation circuit 
 font_test_gen font_gen_unit
 (.clk(clk), video_on(video_on), pixel_x(pixel_x),
  .pixel_y(pixel_y), .rgb_text(rgb_next));
  
  // rgb buffer
  always @(posedge clk)
    if(pixel_tick)
        rgb_reg <= rgb_next;
   // output 
   assign rgb = rgb_reg;
endmodule
