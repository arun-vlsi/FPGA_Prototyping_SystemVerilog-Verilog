`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 13.10.2025 15:23:47
// Design Name: 
// Module Name: dot_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module dot_top
(
input wire clk, reset,
inout wire [1:0] btn,
input wire [2:0] sw,
output wire hsync, vsync,
output wire [2:0] rgb
);

// signal declaration 
wire [9:0] pixel_x, pixel_y;
wire video_on, pixel_tick;
reg [2:0] rgb_reg;
wire [2:0] rgb_next;

// body 
// instantiate VGA sync circuit 
vga_sync vsync_unit 
(.clk(clk), .reset(reset), .hsync(hsync), .vsync(vsync),
 .video_on(video_on), .p_tick(pixel_tick),
 .pixel_x(pixel_x), .pixel_y(pixel_y));
 
 // instantiate graphic generator 
 bitmap_gen bitmap_unit 
   (.clk(clk), .reset(reset), .btn(btn), .sw(sw), 
    .video_on(video_on), .pix_x(pixel_x),
    .pix_y(pixel_y), .bit_rgb(rgb_next));
    
 // rgb buffer
 always @(posedge clk)
   if(pixel_tick)
      rgb_reg <= rgb_next;
  // output 
  assign rgb = rgb_reg;
  
endmodule
