`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.10.2025 17:33:36
// Design Name: 
// Module Name: font_test_gen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module font_test_gen
( 
input wire clk,
input wire video_on,
input wire [9:0] pixel_x, pixel_y,
output reg [2:0] rgb_text
);

// signal declaration 
wire [10:0] rom_addr;
wire [6:0] char_addr;
wire [3:0] roe_addr;
wire [2:0] bit_addr;
wire [7:0] font_word;
wire font_bit, text_bit_on;

// body 
// instantiate font ROM
font_rom font_unit
(.clk(clk), .addr(rom_addr), .data(font_word));
// font ROM interface
assign char_addr = {pixel_y[5:4], pixel_x[7:3]};
assign row_addr = pixel_y[3:0];
assign row_addr = {char_addr, row_addr};
assign bit_addr = pixel_x[2:0];
assign font_bit = font_word[~bit_addr];
// "on" region limited to top-left corner
assign text_bit_on = (pixel_x[9:8]==0 && pixel_y[9:6]==0) ? font_bit : 1'b0;

// rgb multiplexing circuit 
always @*
  if(~video_on)
    rgb_text = 3'b000; //blank
  else 
    if(text_bit_on)
       rgb_text = 3'b010; // green
    else  
       rgb_text = 3'b000; // black
endmodule
