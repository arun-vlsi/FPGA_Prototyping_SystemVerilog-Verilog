`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 16.10.2025 12:24:02
// Design Name: 
// Module Name: text_screen_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module text_screen_top
(
input wire clk, reset,
input wire [2:0] btn,
input wire [6:0] sw,
output wire hsync, vsync,
output wire [2:0] rgb 
);

// signal declaration 
wire [9:0] pixel_x, pixel_y;
wire video_on, pixel_tick;
reg [2:0] rgb_reg;
wire [2:0] rgb_next;
// body 
// instantiate vga sync circuit
vga_sync vsync_unit
(.clk(clk), .reset(reset), .hsync(hsync), .vsync(vsync),
 .video_on(video_on), .p_tick(pixel_tick), 
 .pixel_x(pixel_x), .pixel_y(pixel_y));
 // font generation circuit
 text_screen_gen text_gen_unit
 (.clk(clk), .reset(reset), .video_on(video_on), 
  .btn(btn), .sw(sw), .pixel_x(pixel_x), .pixel_y(pixel_y),
  .text_rgb(rgb_next));
 // rgb buffer
 always @(posedge clk)
    if (pixel_tick)
       rgb_reg <= rgb_next;
 // output 
 assign rgb = rgb_reg;
endmodule
